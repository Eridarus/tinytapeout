module top_level#(
	parameter H_PIXELS = 640,
	parameter V_PIXELS = 480
)
(
	input [3:0] buttons,
	input reset,
	input pix_clk,
	output [1:0] red,
	output [1:0] blu,
	output [1:0] grn,
	output hsync,
	output vsync
);
	
	

endmodule